* File name: C:\Users\user\Desktop\ddd.sch
* Software version: DSCH 2.7a
* Created 04-12-2023 15:30:04
*
* Voltage and current sources
*
V1 3 0 DC 0.6 AC 1 0
V2 4 0 DC 1.2 AC 1 0
vdd 1 0 DC 1.2
*
* Passive devices
*
C1 5 0 0.01nf
*
* Active devices
*
MP1 2 2 1 2 MP W=5u L=0.12u
MN1 2 3 0 2 MN W=5u L=0.12u
MN2 0 4 5 0 MN W=5u L=0.12u
MP2 1 2 5 1 MP W=5u L=0.12u
*
* Warning: "spice.lib" not found, model not declared
.TRAN 0.1ns 250ns
*--WinSpice3--
* Run simulation
*#run
*
* Dump time and volts in "ddd.txt"
*#set nobreak
*#print  V(5)  > ddd.txt
* Show the result in a window
*#plot  V(5) 
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
